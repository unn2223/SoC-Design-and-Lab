`define DATA_WIDTH 8
`define DEPTH_LG2  4
`define REPEAT     20
